`timescale 1ns/1ps

module even_odd_ac;

endmodule
