class instr_coverage extends uvm_subscriber #(instruction);
    `uvm_component_utils(instr_coverage)

    uvm_analysis_imp #(instruction, instr_coverage) imp;
    instruction instr, prev_instr;


    covergroup instr_fields_cg;
        // Opcode
        opcode_cp : coverpoint instr.opcode {
            bins RTYPE = {6'h00};
            bins LW  = {6'h23};
            bins SW  = {6'h2B};
            bins BEQ = {6'h04};
        }

        // Function code
        funct_cp : coverpoint instr.funct {
            bins NOP = {6'h00};
            bins ADD = {6'h20};
            bins AND = {6'h24};
        }

        // ADD
        add_rs : coverpoint instr.rs iff (instr.opcode == 6'h00 && instr.funct == 6'h20) {
            bins rs_vals[] = {[0:4]};
        }
        add_rt : coverpoint instr.rt iff (instr.opcode == 6'h00 && instr.funct == 6'h20) {
            bins rt_vals[] = {[0:4]};
        }
        add_rd : coverpoint instr.rd iff (instr.opcode == 6'h00 && instr.funct == 6'h20) {
            bins rd_vals[] = {[0:4]};
        }
        add_cross : cross add_rs, add_rt, add_rd iff (instr.rd == 5'd0);

        // AND
        and_rs : coverpoint instr.rs iff (instr.opcode == 6'h00 && instr.funct == 6'h24) {
            bins rs_vals[] = {[0:4]};
        }
        and_rt : coverpoint instr.rt iff (instr.opcode == 6'h00 && instr.funct == 6'h24) {
            bins rt_vals[] = {[0:4]};
        }
        and_rd : coverpoint instr.rd iff (instr.opcode == 6'h00 && instr.funct == 6'h24) {
            bins rd_vals[] = {[0:4]};
        }
        and_cross : cross and_rs, and_rt, and_rd iff (instr.rd == 5'd0);

        // LW
        lw_rs : coverpoint instr.rs iff (instr.opcode == 6'h23) {
            bins rs_vals[] = {0};
        }
        lw_rt : coverpoint instr.rt iff (instr.opcode == 6'h23) {
            bins rt_vals[] = {[0:4]};
        }
        lw_imm : coverpoint instr.imm iff (instr.opcode == 6'h23) {
            bins imm_vals[] = {16'h0, 16'h4, 16'h8, 16'hC};
        }
        lw_cross : cross lw_rs, lw_rt, lw_imm;

        // SW
        sw_rs : coverpoint instr.rs iff (instr.opcode == 6'h2B) {
            bins rs_vals[] = {0};
        }
        sw_rt : coverpoint instr.rt iff (instr.opcode == 6'h2B) {
            bins rt_vals[] = {[0:4]};
        }
        sw_imm : coverpoint instr.imm iff (instr.opcode == 6'h2B) {
            bins imm_vals[] = {16'h0, 16'h4, 16'h8, 16'hC};
        }
        sw_cross : cross sw_rs, sw_rt, sw_imm;

        // BEQ
        beq_rs : coverpoint instr.rs iff (instr.opcode == 6'h04) {
            bins rs_vals[] = {[0:4]};
        }
        beq_rt : coverpoint instr.rt iff (instr.opcode == 6'h04) {
            bins rt_vals[] = {[0:4]};
        }
        beq_imm : coverpoint instr.imm iff (instr.opcode == 6'h04) {
            bins imm_vals[] = {16'd1, 16'd2, 16'd3, 16'd4};
        }
        beq_cross : cross beq_rs, beq_rt, beq_imm;
    endgroup


    covergroup branching_cg;
        branch_taken : coverpoint instr.rs {
            bins rs_eq_rt[] = {[0:4]} iff (instr.rs == instr.rt && instr.opcode == 6'h04);
        }
        branch_not_taken_rs : coverpoint instr.rs {
            bins rs_ne_rt[] = {[0:4]} iff (instr.rs != instr.rt && instr.opcode == 6'h04);
        }
        branch_not_taken_rt : coverpoint instr.rt {
            bins rt_ne_rs[] = {[0:4]} iff (instr.rs != instr.rt && instr.opcode == 6'h04);
        }
    endgroup


    covergroup instr_gap_cg;

    function new(string name, uvm_component parent);
        super.new(name, parent);
        $display("Creating instruction coverage collector");
        imp = new("imp", this);
        instr_fields_cg = new();
        branching_cg = new();
    endfunction


    virtual function void write(instruction t);
        instr = t;
        instr_fields_cg.sample();
        branching_cg.sample();
    endfunction
endclass
