module FPAddSub_PrealignModule(
    input  logic [31:0] A,          // Input A, a 32-bit floating point number
    input  logic [31:0] B,          // Input B, a 32-bit floating point number
    input  logic        operation,
    output logic        Sa,         // A's sign
    output logic        Sb,         // B's sign
    output logic [9:0]  ShiftDet,
    output logic [4:0]  InputExc,   // Input numbers are exceptions
    output logic [30:0] Aout,
    output logic [30:0] Bout,
    output logic        Opout
);
	
	// Internal signals
	wire ANaN;			// A is a NaN (Not-a-Number)
	wire BNaN;          // B is a NaN
	wire AInf;			// A is infinity
	wire BInf;			// B is infinity
	wire [7:0] DAB;		// ExpA - ExpB					
	wire [7:0] DBA;     // ExpB - ExpA	
	
	assign ANaN = &(A[30:23]) & |(A[22:0]);		// All one exponent and not all zero mantissa - NaN
	assign BNaN = &(B[30:23]) & |(B[22:0]);		// All one exponent and not all zero mantissa - NaN
	assign AInf = &(A[30:23]) & ~|(A[22:0]);	// All one exponent and all zero mantissa - Infinity
	assign BInf = &(B[30:23]) & ~|(B[22:0]);    // All one exponent and all zero mantissa - Infinity
	
	// Put all flags into exception vector
	assign InputExc = {(ANaN | BNaN | AInf | BInf), ANaN, BNaN, AInf, BInf};
	
	assign DAB = (A[30:23] + ~(B[30:23]) + 1);
	assign DBA = (B[30:23] + ~(A[30:23]) + 1);
	
	assign Sa = A[31];						// A's sign bit
	assign Sb = B[31];						// B's sign	bit
	assign ShiftDet = {DBA[4:0], DAB[4:0]}; // Shift data
	assign Opout = operation;
	assign Aout = A[30:0];
	assign Bout = B[30:0];
	
endmodule
