/*--------------------------------------------------------------
 *  File Name 	: apb_defines.svh
 *  Title 		: This file contains general defines used in APB UVCs 	
 *  Author		: sefaveske@gmail.com	
 *  Date		: 08/24/2018
 *
 *               ##     ####   #    #
 *              #  #   #       #    #
 *             #    #   ####   #    #
 *             ######       #  #    #
 *             #    #  #    #   #  #
 *             #    #   ####     ##
 * ------------------------------------------------------------*/

`ifndef _APB_DEFINES_
`define _APB_DEFINES_

`define ADDR_WIDTH 4                // APB PADDR BUS width           
`define DATA_WIDTH 16               // APB PWDATA and PRDATA Bus width

`endif