module dpi_checker (
    write_if write,     // Push interface
    read_if  read       // Pop interface
);

endmodule
