`timescale 1ns/1ps

module tb_even_odd_ac;

endmodule;
