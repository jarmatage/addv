package memory_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "memory_defines.svh"
    `include "memory_seq_item.svh"
    `include "memory_seq.sv"
    `include "memory_sequencer.svh"
    `include "memory_driver.svh"
    `include "memory_slave_agent.svh"

endpackage