typedef enum {READ, WRITE} mem_agent_mode_t;
