////////////////////////////////////////////////////////////////////////////
// ========================================================================
// This file has the following module implementations:
// 1. top
// 2. mips
// 3. dmem
// 4. imem
// =========================================================================
////////////////////////////////////////////////////////////////////////////
// Top Module 
//  - This module connects the MIPS processor to instruction and data memory
////////////////////////////////////////////////////////////////////////////
module top (
    input clk, reset,
    output [31:0] writedata, dataadr,
    output memwrite
);
    wire [31:0] pc, instr, readdata;

    // instantiate processor and memories
    mips mips (clk, reset, pc, instr, memwrite, dataadr, writedata, readdata);
    imem imem (pc[7:2], instr);
    dmem dmem (clk, memwrite, dataadr, writedata, readdata);
endmodule


//////////////////////////////////////////////////////////////////////
// Single-cycle MIPS Processor Module
//////////////////////////////////////////////////////////////////////
module mips (
    input           clk, reset,
    output  [31:0]  pc,
    input   [31:0]  instr,
    output          memwrite,
    output  [31:0]  aluout, writedata,
    input   [31:0]  readdata
);

    wire memtoreg, branch, alusrc, regdst, regwrite, jump;
    wire [2:0] alucontrol;

    controller c(instr[31:26], instr[5:0], zero, memtoreg, memwrite, pcsrc, alusrc, regdst, regwrite, jump, alucontrol);

    datapath dp(clk, reset, memtoreg, pcsrc, alusrc, regdst, regwrite, jump,alucontrol, zero, pc, instr, aluout, writedata, readdata);
endmodule


//////////////////////////////////////////////////////////////////////
// Data Memory Module
// - Uses 32x64 SRAM model generated by OpenRAM 
//////////////////////////////////////////////////////////////////////
module dmem (
    input clk, we,
    input [31:0] a, wd,
    output [31:0] rd
);
    // OpenRAM signals
    wire csb0;          // Chip select (active low)
    wire web0;          // Write enable (active low)
    wire [5:0] addr0;   // 6-bit address
    wire [31:0] din0;   // Data input
    wire [31:0] dout0;  // Data output
    

    assign csb0 = 1'b0;         // Always enabled
    assign web0 = ~we;          // Invert we (active high to active low)
    assign addr0 = a[7:2];      // Word-aligned address (6 bits)
    assign din0 = wd;           // Write data
    assign rd = dout0;          // Read data
    
    // OpenRAM instantiation
    SRAM_32x64_1rw dmem_ram (
        .clk0(clk),
        .csb0(csb0),
        .web0(web0),
        .addr0(addr0),
        .din0(din0),
        .dout0(dout0)
    );
endmodule


//////////////////////////////////////////////////////////////////////
// Instruction Memory Module
// - Uses 32x64 SRAM model generated by OpenRAM 
//////////////////////////////////////////////////////////////////////
module imem (
    input [5:0] a,
    output [31:0] rd
);
    // OpenRAM interface signals
    wire clk0;          // Clock
    wire csb0;          // Chip select (active low)
    wire web0;          // Write enable (active low)
    wire [5:0] addr0;   // 6-bit address
    wire [31:0] din0;   // Data input
    wire [31:0] dout0;  // Data output
    
    // Control signal connections
    assign clk0 = 1'b0;         // No clock needed for read-only
    assign csb0 = 1'b0;         // Always enabled
    assign web0 = 1'b1;         // Always read (never write)
    assign addr0 = a;           // Address from processor
    assign din0 = 32'b0;        // No data to write
    assign rd = dout0;          // Read data
    
    // OpenRAM instantiation
    SRAM_32x64_1rw imem_ram (
        .clk0(clk0),
        .csb0(csb0),
        .web0(web0),
        .addr0(addr0),
        .din0(din0),
        .dout0(dout0)
    );
endmodule