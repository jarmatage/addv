typedef enum {READ, WRITE} mem_agent_mode_t;
typedef bit [31:0] mem_array_t[*];
