class serialalu_configuration extends uvm_object;
	`uvm_object_utils(serialalu_configuration)

	function new(string name = "");
		super.new(name);
	endfunction: new
endclass: serialalu_configuration
